////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module      : top.sv
// Project      : M.Tech-VLSI-Main-Project-Adder_Verification
// Description: 
// This is the top module.
// It connects the DUT and testbench.
// Firstly, the interface is instantiated with the clk and reset signals.
// Then, the interface is passed as a parameter to the program block.
// And lastly, the DUT is invoked with port declarations made with respect to interface signals.
//
// Change history: 18/05/20 - V1.0 Initial working version created  (owner: Abhishek Kumar)
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module top;
	bit clk, reset;

	always #5 clk = ~clk;

	intf_adr intf_1(clk, reset);
	test test_1(intf_1);
	adder DUT (
	  .clk (intf_1.clk),
	  .reset (intf_1.reset),
	  .a (intf_1.a),
	  .b (intf_1.b),
	  .c (intf_1.c)
	  );
	  
	initial begin
	reset = 1 ; clk = 0; 
	#30; reset = 0;
	end
	  
	initial
	begin
	$dumpfile ("dump.vcd");
	$dumpvars;
	end

endmodule