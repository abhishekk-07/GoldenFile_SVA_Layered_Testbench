////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module      : interface.sv
// Project      : M.Tech-VLSI-Main-Project-Adder_Verification
// Description: 
// This is the interface module.
// Two signals are taken as input for the interface, clk and reset.
// Rest of the signals are mentioned as logic.
// For the purpose of measuring the coverage, there is a covergroup, cg, defined in the interface for all the variables.
//
// Change history: 18/05/20 - V1.0 Initial working version created  (owner: Abhishek Kumar)
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

interface intf_adr( input logic clk, reset);
  logic [3:0] a;
  logic [3:0] b;
  logic [4:0] c;
  
  covergroup cg @ (posedge clk);
    cov_a : coverpoint a;
    cov_b : coverpoint b;
    cov_c : coverpoint c;
  endgroup 
  
  cg cg_1 = new();
  
  
endinterface
