////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module      : monitor.sv
// Project      : M.Tech-VLSI-Main-Project-Adder_Verification
// Description: 
// This is the monitor module.
// It transmits a sampled interface signal to the scoreboard via the mailbox (mon2scb).
// The constructor takes two parameters, a virtual interface and a mailbox handle.
//
// Change history: 18/05/20 - V1.0 Initial working version created  (owner: Abhishek Kumar)
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`include "driver.sv"
class monitor;
   virtual intf_adr vif;
   mailbox mon2scb;
   
   function new ( virtual intf_adr vif, mailbox mon2scb);
     this.vif = vif;
     this.mon2scb = mon2scb;
   endfunction
   
   task main;
     forever
     begin
       transaction trans;
       trans = new();
       @ (posedge vif.clk)
       trans.a = vif.a;
       trans.b = vif.b;
       trans.c = vif.c;
       mon2scb.put(trans);
     end
   endtask
   
 endclass