////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Module      : transaction.sv
// Project      : M.Tech-VLSI-Main-Project-Adder_Verification
// Description: 
// This is the transactor module. 
// It provides randomized inputs to the design.
// There are two inputs and one output declared in this module.
// Inputs are a and b.
// Output is c.
//
// Change history: 18/05/20 - V1.0 Initial working version created  (owner: Abhishek Kumar)
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class transaction;
  randc bit [3:0] a;
  rand bit [3:0] b;
          bit [4:0] c;
endclass